module main
import argile

fn main() {
	println('Hello World!')
	println(argile.clay__max(5.2, 10))
	println(argile.clay__min(5.2, 10))
}