module argile

